

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity MUL8bit is
end MUL8bit;

--}} End of automatically maintained section

architecture MUL8bit of MUL8bit is
begin

	 -- enter your statements here --

end MUL8bit;
